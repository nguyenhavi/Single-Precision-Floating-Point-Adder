`timescale 1ns / 1ps
module FloatingPointAdder_tb;

reg [31:0] A;
reg [31:0] B;

wire [31:0] Out;

FloatingPointAdder uut (.A(A), .B(B), .Out(Out));

initial begin

	A = 32'b01000001001101100000000000000001;//11.375
	B = 32'b01000000101100100000010000011011;//5.56300
	//SUM = 16.938
	
	// Wait 200 ns to new state
	#200
	A = 32'b01000000101110000000000000000000; // 5.75
	B = 32'b01000000010100000000000000000000; // 3.25
	//SUM = 9
	#200 
	A=32'b01000010011011111110101110000101;//59.979
	B=32'b01000000110100000000000000000000;//6.5
	//SUM = 66.479
		 
	#200 
	A=32'b01000100011110100010000000000000;//1000.5
	B=32'b01000100011101010110100111011011;//981.654
	//SUM = 1982.1539
		 
	#200
	A=32'b01000100000010010111111100101011;//549.987
	B=32'b01000000101100100000010000011001;//5.563
	//SUM = 555.499
		
end
      
endmodule

